LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY reg IS
   PORT(
			A        : IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
			res, clk : IN  STD_LOGIC;
			Q        : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
   );
END reg;

ARCHITECTURE behavior OF reg IS
BEGIN

	PROCESS(res, clk)
   BEGIN
		IF res = '0' THEN
			Q <= "00000000";
      ELSIF(clk'EVENT AND clk = '1') THEN
			Q <= A;
		END IF;
   END PROCESS;
	
END behavior;